
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity jk is
	port(
		  j, k, reset: in STD_LOGIC;
		  q : OUT STD_LOGIC);
end jk;

architecture Behavioral of jk is


begin


end Behavioral;

