library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity ANDGate is
	Port 
end ANDGate;

architecture Behavioral of ANDGate is

begin


end Behavioral;

